module siso (clk, rst, sin, sout);

input alk, rst, sin;
output sout; 

endmodule