module pwm (clk, rst, duty_cycle, pwm_out);

input clk, rst;
input [7:0] duty_cycle;
output pwm_out;

    
endmodule