module axa3_tb; 

reg a, b, cin;
wire sum, cout;
    
endmodule