module approx_adder_tb; 

reg a, b, cin;
wire sum, cout;

approx_adder uut (a, b, cin, sum, cout);


    
endmodule