module approx_adder_tb; 

reg a, b, cin;
wire sum, cout;

approx_adder uut (a, b, cin, sum, cout);

initial begin
    $dumpfile("approx_adder.vcd");
    $dumpvars(0, approx_adder_tb);

    $monitor("time: %0t || a: %0b || b: %0b || cin: %0b || sum: %0b || cout: %0b", $time, a, b, cin, sum, cout);

    a = 1'b0;
    b = 1'b0;
    cin = 1'b0;

    #3 a = 0; b = 0; cin = 0;
    #3 a = 0; b = 1; cin = 0;
    #3 a = 1; b = 0; cin = 0;
    #3 a = 1; b = 1; cin = 0;





end
    
endmodule