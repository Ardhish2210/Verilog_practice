module pulse (clk, rst, in_pulse, out_pulse);

input clk, rst, in_pulse;
output out_pulse;

    
endmodule