$date
	Sun Aug 24 17:04:28 2025
$end
$version
	Icarus Verilog
$end
$timescale
	1ns
$end
$scope module xor_using_nand_tb $end
$var wire 1 ! y $end
$var reg 1 " a $end
$var reg 1 # b $end
$upscope $end
$enddefinitions $end
$comment Show the parameter values. $end
$dumpall
$end
#0
$dumpvars
0#
0"
z!
$end
#10
1#
#20
0#
1"
#30
1#
#40
