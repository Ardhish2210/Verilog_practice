module ama2 (a, b, cin, sum, cout);

input a, b, cin;
output sum, cout;


    
endmodule