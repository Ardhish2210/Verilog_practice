module counter_ten (clk, rst, counter);

input clk, rst;
output counter;

    
endmodule