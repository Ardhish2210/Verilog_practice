module priority_encoder_new (d, out, valid);
    
input valid;
input [7:0] d;
output [2:0] out;


endmodule