module ama4 #(
    parameters
) (
    ports
);
    
endmodule