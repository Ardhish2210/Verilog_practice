module approx_adder_tb; 

reg a, b, cin;
wire sum, cout;
    
endmodule