module encoder (a, enable, out);

input [2:0] a;
input enable;
output [7:0] out;

always@(*) begin
    
end
    
endmodule