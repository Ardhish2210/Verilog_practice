module (sel, enable, a, bus_line);

input [1:0] sel;
input enable;
input [3:0] a;
output bus_line;

endmodule