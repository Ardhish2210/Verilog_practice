module approx_adder (a, b, cin, sum, cout);
    
endmodule