module mood #(
    parameters
) (
    ports
);
    
endmodule