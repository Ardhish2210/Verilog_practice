module counter_ten ();
    
endmodule