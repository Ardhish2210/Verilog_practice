module ripple_carry_two (a, b, cin, sum, cout);

input 
    
endmodule