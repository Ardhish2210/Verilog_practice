module ripple_adder (a, b, cin, sum, cout);

input cin;
input [3:0] a, b;
output sum, cout;

    
endmodule