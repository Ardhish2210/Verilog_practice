module full_adder #(
    parameters
) (
    ports
);
    
endmodule