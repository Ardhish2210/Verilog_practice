module counter_ten (clk, rst, counter);

input clk, rst;
output counter;

always @(posedge clk or posedge rst) begin
    if(rst) begin
        
    end

end


    
endmodule