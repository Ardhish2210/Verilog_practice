module cla (a, b, sum, cout);

input [3:0] a, b;
output [3:0] sum;
wire [3:0] P, G; // P = propagation carry, G = Generated carry




endmodule