module full_adder(a, b, cin, sum, cout);

// In this module I will make the full adder cicuit using the gate level modeling (structural modeling)

input a, b, cin;
output sum, cout;

endmodule