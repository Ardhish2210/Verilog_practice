`timescale 1ns/1ns
`include "pwm.v"

module pwm_tb;

reg clk, rst;
reg [7:0] duty_cycle;
wire pwm_out;
    
endmodule