module esa3 (a, b, sum);

input [7:0] a, b;
output [8:0] sum;


    
endmodule