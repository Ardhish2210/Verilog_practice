module axa3_tb; 

reg a, b, cin;
wire sum, cout;

axa3 uut (a, b, cin, sum, cout);

    
endmodule