module esa3_tb; 

reg [7:0] a,b;
wire [8:0] sum;

endmodule