`timescale 1ns/1ns
`include "encoder.v"

module encoder_tb; 

reg [2:0] a;
reg enable;
wire [7:0] out;

encoder uut (a, enable, out);

initial begin

    $dumpfile("encoder.vcd");
    $dumpvars(0, encoder_tb);

    $monitor("Time: %0t || a: %b || enable: %b || out: %b", $time, a, enable, out);

    a = 3'b000; enable = 0;
    
    #5 a = 3'b010; enable = 1;
    #5 a = 3'b110; enable = 1;
    #5 a = 3'b011; enable = 1;
    #5 a = 3'b101; enable = 1;

    #10 $finish;
end
    
endmodule