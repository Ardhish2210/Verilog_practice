module new_adder (a, b, sum);

input [31:0] a, b;
output [32:0] sum;
    
endmodule