module eta6_tb;

reg [5:0] A, B;
wire [5:0] SUM;
wire COUT;

    
endmodule