`timescale 1ns/1ns
`include "xor_using_nand.v"

module xor_using_nand_tb;

reg a, b;
wire y;


endmodule