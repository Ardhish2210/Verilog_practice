module xor_using_nand (a, b, y);

input a, b;
output y;

wire d, e, f;

endmodule