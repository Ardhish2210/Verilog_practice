module one_hot_encoder_tb;

reg [3:0]
endmodule