module eta6 (A, B, SUM, COUT);

input [5:0] A, B;
output [5:0] SUM;
output COUT;

     
endmodule