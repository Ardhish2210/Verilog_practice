module majority_gate (a, b, c, out);

input a, b, c;
output out;

//This is basically like VOTING MACHINE, The output will be 1 if there are majority 1's in the input and 0 if there are majority 0's in the input
endmodule