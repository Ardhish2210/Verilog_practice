module(a, out);

input [3:0] a;
output [7:0] out;



endmodule