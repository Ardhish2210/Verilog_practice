module mood_tb; 


mood uut (brain_wave, clk, rst, rgb, blink);


    
endmodule