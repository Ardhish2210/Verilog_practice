module carry_save_adder #(
    parameters
) (
    ports
);
    
endmodule