`timescale 1ns/1ns
`include "ama2.v"

module ama2_tb; 

reg a, b, cin;
wire sum, cout;

    
endmodule