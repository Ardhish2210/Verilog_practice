module xor_using_nand (a, b, y);


endmodule