module majority_gate (a, b, c, out);

input a, b, c;
output out;

endmodule