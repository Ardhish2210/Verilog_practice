`timescale 1ns/1ns
`include "counter_ten.v"

module counter_ten_tb; 

reg clk, rst;
wire [3:0] counter;

endmodule